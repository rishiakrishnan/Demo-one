file_input("output","DebugSoc","DebugSoc","bsv")
file_input("output","mixed_cluster","mixed_cluster","bsv")
file_input("output","pinmux_axi4lite","pinmux_axi4lite","bsv")
file_input("output","pinmux","pinmux","bsv")
file_input("output","pwm_cluster","pwm_cluster","bsv")
file_input("output","sign_dump","sign_dump","bsv")
file_input("output","Soc","Soc","bsv")
file_input("output","spi_cluster","spi_cluster","bsv")
file_input("output","TbSoc","TbSoc","bsv")
file_input("output","uart_cluster","uart_cluster","bsv")
file_input("output","dsoc","Soc","defines")