
/*
   This BSV file has been generated by the PinMux tool available at:
   https://bitbucket.org/casl/pinmux.

   Authors: Neel Gala, Luke
   Date of generation: Fri Aug 23 12:07:59 2024
*/

package pinmux;

   typedef struct{
      Bit#(1) outputval;      // output from core to pad                bit7
      Bit#(1) output_en;      // output enable from core to pad         bit6
      Bit#(1) input_en;       // input enable from core to io_cell      bit5
      Bit#(1) pullup_en;      // pullup enable from core to io_cell     bit4
      Bit#(1) pulldown_en;    // pulldown enable from core to io_cell   bit3
      Bit#(1) drivestrength;  // drivestrength from core to io_cell     bit2
      Bit#(1) pushpull_en;    // pushpull enable from core to io_cell   bit1
      Bit#(1) opendrain_en;   // opendrain enable form core to io_cell  bit0
   } GenericIOType deriving(Eq,Bits,FShow);

   interface MuxSelectionLines;

      // declare the method which will capture the user pin-mux
      // selection values.The width of the input is dependent on the number
      // of muxes happening per IO. For now we have a generalized width
      // where each IO will have the same number of muxes.
     method  Action cell0_mux (Bit#(2) in);
     method  Action cell1_mux (Bit#(2) in);
     method  Action cell2_mux (Bit#(1) in);
     method  Action cell3_mux (Bit#(1) in);
     method  Action cell8_mux (Bit#(1) in);
     method  Action cell9_mux (Bit#(1) in);
     method  Action cell10_mux (Bit#(1) in);
     method  Action cell11_mux (Bit#(1) in);
     method  Action cell12_mux (Bit#(1) in);
     method  Action cell13_mux (Bit#(1) in);
      endinterface

      interface PeripheralSide;
      // declare the interface to the IO cells.
      // Each IO cell will have 8 input field (output from pin mux
      // and on output field (input to pinmux)
          // interface declaration between IO-0 and pinmux
    (*always_ready*) method  GenericIOType io0_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io0_inputval (Bit#(1) in);
          // interface declaration between IO-1 and pinmux
    (*always_ready*) method  GenericIOType io1_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io1_inputval (Bit#(1) in);
          // interface declaration between IO-2 and pinmux
    (*always_ready*) method  GenericIOType io2_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io2_inputval (Bit#(1) in);
          // interface declaration between IO-3 and pinmux
    (*always_ready*) method  GenericIOType io3_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io3_inputval (Bit#(1) in);
          // interface declaration between IO-4 and pinmux
    (*always_ready*) method  GenericIOType io4_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io4_inputval (Bit#(1) in);
          // interface declaration between IO-5 and pinmux
    (*always_ready*) method  GenericIOType io5_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io5_inputval (Bit#(1) in);
          // interface declaration between IO-6 and pinmux
    (*always_ready*) method  GenericIOType io6_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io6_inputval (Bit#(1) in);
          // interface declaration between IO-7 and pinmux
    (*always_ready*) method  GenericIOType io7_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io7_inputval (Bit#(1) in);
          // interface declaration between IO-8 and pinmux
    (*always_ready*) method  GenericIOType io8_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io8_inputval (Bit#(1) in);
          // interface declaration between IO-9 and pinmux
    (*always_ready*) method  GenericIOType io9_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io9_inputval (Bit#(1) in);
          // interface declaration between IO-10 and pinmux
    (*always_ready*) method  GenericIOType io10_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io10_inputval (Bit#(1) in);
          // interface declaration between IO-11 and pinmux
    (*always_ready*) method  GenericIOType io11_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io11_inputval (Bit#(1) in);
          // interface declaration between IO-12 and pinmux
    (*always_ready*) method  GenericIOType io12_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io12_inputval (Bit#(1) in);
          // interface declaration between IO-13 and pinmux
    (*always_ready*) method  GenericIOType io13_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io13_inputval (Bit#(1) in);
          // interface declaration between IO-14 and pinmux
    (*always_ready*) method  GenericIOType io14_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io14_inputval (Bit#(1) in);
          // interface declaration between IO-15 and pinmux
    (*always_ready*) method  GenericIOType io15_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io15_inputval (Bit#(1) in);
          // interface declaration between IO-16 and pinmux
    (*always_ready*) method  GenericIOType io16_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io16_inputval (Bit#(1) in);
          // interface declaration between IO-17 and pinmux
    (*always_ready*) method  GenericIOType io17_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io17_inputval (Bit#(1) in);
          // interface declaration between IO-18 and pinmux
    (*always_ready*) method  GenericIOType io18_cell;
    (*always_ready,always_enabled,result="io"*) method 
                       Action io18_inputval (Bit#(1) in);
          // interface declaration between UART-0 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) uart0_rx;
    (*always_ready,always_enabled*) method  Action uart0_tx (Bit#(1) in);
          // interface declaration between UART-1 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) uart1_rx;
    (*always_ready,always_enabled*) method  Action uart1_tx (Bit#(1) in);
          // interface declaration between UART-2 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) uart2_rx;
    (*always_ready,always_enabled*) method  Action uart2_tx (Bit#(1) in);
          // interface declaration between UART-3 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) uart3_rx;
    (*always_ready,always_enabled*) method  Action uart3_tx (Bit#(1) in);
          // interface declaration between SPI-0 and pinmux
    (*always_ready,always_enabled*) method  Action spi_sclk (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action spi_mosi (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action spi_ss (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) spi_miso;
          // interface declaration between TWI-0 and pinmux
    (*always_ready,always_enabled*) method  Action twi0_sda_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action twi0_sda_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) twi0_sda_in;
    (*always_ready,always_enabled*) method  Action twi0_scl_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action twi0_scl_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) twi0_scl_in;
          // interface declaration between TWI-1 and pinmux
    (*always_ready,always_enabled*) method  Action twi1_sda_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action twi1_sda_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) twi1_sda_in;
    (*always_ready,always_enabled*) method  Action twi1_scl_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action twi1_scl_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) twi1_scl_in;
          // interface declaration between SD-0 and pinmux
    (*always_ready,always_enabled*) method  Action sd0_clk (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_cmd (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_d0_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_d0_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd0_d0_in;
    (*always_ready,always_enabled*) method  Action sd0_d1_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_d1_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd0_d1_in;
    (*always_ready,always_enabled*) method  Action sd0_d2_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_d2_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd0_d2_in;
    (*always_ready,always_enabled*) method  Action sd0_d3_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd0_d3_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd0_d3_in;
          // interface declaration between SD-1 and pinmux
    (*always_ready,always_enabled*) method  Action sd1_clk (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_cmd (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_d0_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_d0_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd1_d0_in;
    (*always_ready,always_enabled*) method  Action sd1_d1_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_d1_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd1_d1_in;
    (*always_ready,always_enabled*) method  Action sd1_d2_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_d2_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd1_d2_in;
    (*always_ready,always_enabled*) method  Action sd1_d3_out (Bit#(1) in);
    (*always_ready,always_enabled*) method  Action sd1_d3_outen (Bit#(1) in);
    (*always_ready,always_enabled*) method  Bit#(1) sd1_d3_in;
          // interface declaration between JTAG-0 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) jtag0_tdi;
    (*always_ready,always_enabled*) method  Bit#(1) jtag0_tms;
    (*always_ready,always_enabled*) method  Bit#(1) jtag0_tclk;
    (*always_ready,always_enabled*) method  Bit#(1) jtag0_trst;
    (*always_ready,always_enabled*) method  Action jtag0_tdo (Bit#(1) in);
          // interface declaration between JTAG-1 and pinmux
    (*always_ready,always_enabled*) method  Bit#(1) jtag1_tdi;
    (*always_ready,always_enabled*) method  Bit#(1) jtag1_tms;
    (*always_ready,always_enabled*) method  Bit#(1) jtag1_tclk;
    (*always_ready,always_enabled*) method  Bit#(1) jtag1_trst;
    (*always_ready,always_enabled*) method  Action jtag1_tdo (Bit#(1) in);
          // interface declaration between PWM-0 and pinmux
    (*always_ready,always_enabled*) method  Action pwm_pwm (Bit#(1) in);
   endinterface

   interface Ifc_pinmux;
      interface MuxSelectionLines mux_lines;
      interface PeripheralSide peripheral_side;
   endinterface
   (*synthesize*)
   module mkpinmux(Ifc_pinmux);

      // the followins wires capture the pin-mux selection
      // values for each mux assigned to a CELL

      Wire#(Bit#(2)) wrcell0_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell1_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell2_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell3_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell8_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell9_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell10_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell11_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell12_mux<-mkDWire(0);
      Wire#(Bit#(2)) wrcell13_mux<-mkDWire(0);
      // following wires capture signals to IO CELL if io-0 is
      // allotted to it
      GenericIOType cell0_mux_out=unpack(0);
      Wire#(Bit#(1)) cell0_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-1 is
      // allotted to it
      GenericIOType cell1_mux_out=unpack(0);
      Wire#(Bit#(1)) cell1_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-2 is
      // allotted to it
      GenericIOType cell2_mux_out=unpack(0);
      Wire#(Bit#(1)) cell2_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-3 is
      // allotted to it
      GenericIOType cell3_mux_out=unpack(0);
      Wire#(Bit#(1)) cell3_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-4 is
      // allotted to it
      GenericIOType cell4_mux_out=unpack(0);
      Wire#(Bit#(1)) cell4_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-5 is
      // allotted to it
      GenericIOType cell5_mux_out=unpack(0);
      Wire#(Bit#(1)) cell5_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-6 is
      // allotted to it
      GenericIOType cell6_mux_out=unpack(0);
      Wire#(Bit#(1)) cell6_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-7 is
      // allotted to it
      GenericIOType cell7_mux_out=unpack(0);
      Wire#(Bit#(1)) cell7_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-8 is
      // allotted to it
      GenericIOType cell8_mux_out=unpack(0);
      Wire#(Bit#(1)) cell8_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-9 is
      // allotted to it
      GenericIOType cell9_mux_out=unpack(0);
      Wire#(Bit#(1)) cell9_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-10 is
      // allotted to it
      GenericIOType cell10_mux_out=unpack(0);
      Wire#(Bit#(1)) cell10_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-11 is
      // allotted to it
      GenericIOType cell11_mux_out=unpack(0);
      Wire#(Bit#(1)) cell11_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-12 is
      // allotted to it
      GenericIOType cell12_mux_out=unpack(0);
      Wire#(Bit#(1)) cell12_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-13 is
      // allotted to it
      GenericIOType cell13_mux_out=unpack(0);
      Wire#(Bit#(1)) cell13_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-14 is
      // allotted to it
      GenericIOType cell14_mux_out=unpack(0);
      Wire#(Bit#(1)) cell14_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-15 is
      // allotted to it
      GenericIOType cell15_mux_out=unpack(0);
      Wire#(Bit#(1)) cell15_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-16 is
      // allotted to it
      GenericIOType cell16_mux_out=unpack(0);
      Wire#(Bit#(1)) cell16_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-17 is
      // allotted to it
      GenericIOType cell17_mux_out=unpack(0);
      Wire#(Bit#(1)) cell17_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if io-18 is
      // allotted to it
      GenericIOType cell18_mux_out=unpack(0);
      Wire#(Bit#(1)) cell18_mux_in<-mkDWire(0);

      // following wires capture signals to IO CELL if uart-0 is
      // allotted to it
      Wire#(Bit#(1)) wruart0_rx<-mkDWire(0);
      Wire#(Bit#(1)) wruart0_tx<-mkDWire(0);
      GenericIOType uart0_rx_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType uart0_tx_io = GenericIOType{
                 outputval:wruart0_tx,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if uart-1 is
      // allotted to it
      Wire#(Bit#(1)) wruart1_rx<-mkDWire(0);
      Wire#(Bit#(1)) wruart1_tx<-mkDWire(0);
      GenericIOType uart1_rx_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType uart1_tx_io = GenericIOType{
                 outputval:wruart1_tx,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if uart-2 is
      // allotted to it
      Wire#(Bit#(1)) wruart2_rx<-mkDWire(0);
      Wire#(Bit#(1)) wruart2_tx<-mkDWire(0);
      GenericIOType uart2_rx_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType uart2_tx_io = GenericIOType{
                 outputval:wruart2_tx,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if uart-3 is
      // allotted to it
      Wire#(Bit#(1)) wruart3_rx<-mkDWire(0);
      Wire#(Bit#(1)) wruart3_tx<-mkDWire(0);
      GenericIOType uart3_rx_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType uart3_tx_io = GenericIOType{
                 outputval:wruart3_tx,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if spi-0 is
      // allotted to it
      Wire#(Bit#(1)) wrspi_sclk<-mkDWire(0);
      Wire#(Bit#(1)) wrspi_mosi<-mkDWire(0);
      Wire#(Bit#(1)) wrspi_ss<-mkDWire(0);
      Wire#(Bit#(1)) wrspi_miso<-mkDWire(0);
      GenericIOType spi_sclk_io = GenericIOType{
                 outputval:wrspi_sclk,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType spi_mosi_io = GenericIOType{
                 outputval:wrspi_mosi,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType spi_ss_io = GenericIOType{
                 outputval:wrspi_ss,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType spi_miso_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if twi-0 is
      // allotted to it
      Wire#(Bit#(1)) wrtwi0_sda_out<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi0_sda_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi0_sda_in<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi0_scl_out<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi0_scl_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi0_scl_in<-mkDWire(0);
      GenericIOType twi0_sda_io = GenericIOType{
                 outputval:wrtwi0_sda_out,
                 output_en:wrtwi0_sda_outen,
                 input_en:~wrtwi0_sda_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType twi0_scl_io = GenericIOType{
                 outputval:wrtwi0_scl_out,
                 output_en:wrtwi0_scl_outen,
                 input_en:~wrtwi0_scl_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if twi-1 is
      // allotted to it
      Wire#(Bit#(1)) wrtwi1_sda_out<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi1_sda_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi1_sda_in<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi1_scl_out<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi1_scl_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrtwi1_scl_in<-mkDWire(0);
      GenericIOType twi1_sda_io = GenericIOType{
                 outputval:wrtwi1_sda_out,
                 output_en:wrtwi1_sda_outen,
                 input_en:~wrtwi1_sda_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType twi1_scl_io = GenericIOType{
                 outputval:wrtwi1_scl_out,
                 output_en:wrtwi1_scl_outen,
                 input_en:~wrtwi1_scl_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if sd-0 is
      // allotted to it
      Wire#(Bit#(1)) wrsd0_clk<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_cmd<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d0_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d0_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d0_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d1_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d1_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d1_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d2_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d2_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d2_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d3_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d3_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd0_d3_in<-mkDWire(0);
      GenericIOType sd0_clk_io = GenericIOType{
                 outputval:wrsd0_clk,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd0_cmd_io = GenericIOType{
                 outputval:wrsd0_cmd,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd0_d0_io = GenericIOType{
                 outputval:wrsd0_d0_out,
                 output_en:wrsd0_d0_outen,
                 input_en:~wrsd0_d0_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd0_d1_io = GenericIOType{
                 outputval:wrsd0_d1_out,
                 output_en:wrsd0_d1_outen,
                 input_en:~wrsd0_d1_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd0_d2_io = GenericIOType{
                 outputval:wrsd0_d2_out,
                 output_en:wrsd0_d2_outen,
                 input_en:~wrsd0_d2_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd0_d3_io = GenericIOType{
                 outputval:wrsd0_d3_out,
                 output_en:wrsd0_d3_outen,
                 input_en:~wrsd0_d3_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if sd-1 is
      // allotted to it
      Wire#(Bit#(1)) wrsd1_clk<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_cmd<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d0_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d0_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d0_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d1_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d1_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d1_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d2_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d2_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d2_in<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d3_out<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d3_outen<-mkDWire(0);
      Wire#(Bit#(1)) wrsd1_d3_in<-mkDWire(0);
      GenericIOType sd1_clk_io = GenericIOType{
                 outputval:wrsd1_clk,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd1_cmd_io = GenericIOType{
                 outputval:wrsd1_cmd,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd1_d0_io = GenericIOType{
                 outputval:wrsd1_d0_out,
                 output_en:wrsd1_d0_outen,
                 input_en:~wrsd1_d0_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd1_d1_io = GenericIOType{
                 outputval:wrsd1_d1_out,
                 output_en:wrsd1_d1_outen,
                 input_en:~wrsd1_d1_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd1_d2_io = GenericIOType{
                 outputval:wrsd1_d2_out,
                 output_en:wrsd1_d2_outen,
                 input_en:~wrsd1_d2_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType sd1_d3_io = GenericIOType{
                 outputval:wrsd1_d3_out,
                 output_en:wrsd1_d3_outen,
                 input_en:~wrsd1_d3_outen,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if jtag-0 is
      // allotted to it
      Wire#(Bit#(1)) wrjtag0_tdi<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag0_tms<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag0_tclk<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag0_trst<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag0_tdo<-mkDWire(0);
      GenericIOType jtag0_tdi_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag0_tms_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag0_tclk_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag0_trst_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag0_tdo_io = GenericIOType{
                 outputval:wrjtag0_tdo,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if jtag-1 is
      // allotted to it
      Wire#(Bit#(1)) wrjtag1_tdi<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag1_tms<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag1_tclk<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag1_trst<-mkDWire(0);
      Wire#(Bit#(1)) wrjtag1_tdo<-mkDWire(0);
      GenericIOType jtag1_tdi_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag1_tms_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag1_tclk_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag1_trst_io = GenericIOType{
                 outputval:0,
                 output_en:0,
                 input_en:1,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };
      GenericIOType jtag1_tdo_io = GenericIOType{
                 outputval:wrjtag1_tdo,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };

      // following wires capture signals to IO CELL if pwm-0 is
      // allotted to it
      Wire#(Bit#(1)) wrpwm_pwm<-mkDWire(0);
      GenericIOType pwm_pwm_io = GenericIOType{
                 outputval:wrpwm_pwm,
                 output_en:1,
                 input_en:0,
                 pullup_en:0,
                 pulldown_en:0,
                 pushpull_en:0,
                 drivestrength:0,
                 opendrain_en:0
      };


      /*====== This where the muxing starts for each io-cell======*/
       cell0_mux_out=wrcell0_mux==0?uart0_tx_io:
			wrcell0_mux==1?spi0_sclk_io:
			wrcell0_mux==2?uart2_tx_io:
			uart3_tx_io;
      cell1_mux_out=wrcell1_mux==0?uart0_rx_io:
			wrcell1_mux==1?spi0_mosi_io:
			wrcell1_mux==2?uart2_rx_io:
			uart3_rx_io;

      rule assign_wruart0_rx_on_cell1(wrcell1_mux==0);
        wruart0_rx<=cell1_mux_in;
      endrule


      rule assign_wruart2_rx_on_cell1(wrcell1_mux==2);
        wruart2_rx<=cell1_mux_in;
      endrule


      rule assign_wruart3_rx_on_cell1(wrcell1_mux==3);
        wruart3_rx<=cell1_mux_in;
      endrule

      cell2_mux_out=wrcell2_mux==0?twi0_sda_io:
			spi0_ss_io;

      rule assign_wrtwi0_sda_in_on_cell2(wrcell2_mux==0);
        wrtwi0_sda_in<=cell2_mux_in;
      endrule

      cell3_mux_out=wrcell3_mux==0?twi0_scl_io:
			spi0_miso_io;

      rule assign_wrtwi0_scl_in_on_cell3(wrcell3_mux==0);
        wrtwi0_scl_in<=cell3_mux_in;
      endrule


      rule assign_wrspi0_miso_on_cell3(wrcell3_mux==1);
        wrspi0_miso<=cell3_mux_in;
      endrule

      cell8_mux_out=wrcell8_mux==0?sd0_clk_io:
			sd1_clk_io;
      cell9_mux_out=wrcell9_mux==0?sd0_cmd_io:
			sd1_cmd_io;
      cell10_mux_out=wrcell10_mux==0?sd0_d0_io:
			sd1_d0_io;

      rule assign_wrsd0_d0_in_on_cell10(wrcell10_mux==0);
        wrsd0_d0_in<=cell10_mux_in;
      endrule


      rule assign_wrsd1_d0_in_on_cell10(wrcell10_mux==1);
        wrsd1_d0_in<=cell10_mux_in;
      endrule

      cell11_mux_out=wrcell11_mux==0?sd0_d1_io:
			sd1_d1_io;

      rule assign_wrsd0_d1_in_on_cell11(wrcell11_mux==0);
        wrsd0_d1_in<=cell11_mux_in;
      endrule


      rule assign_wrsd1_d1_in_on_cell11(wrcell11_mux==1);
        wrsd1_d1_in<=cell11_mux_in;
      endrule

      cell12_mux_out=wrcell12_mux==0?sd0_d2_io:
			sd1_d2_io;

      rule assign_wrsd0_d2_in_on_cell12(wrcell12_mux==0);
        wrsd0_d2_in<=cell12_mux_in;
      endrule


      rule assign_wrsd1_d2_in_on_cell12(wrcell12_mux==1);
        wrsd1_d2_in<=cell12_mux_in;
      endrule

      cell13_mux_out=wrcell13_mux==0?sd0_d3_io:
			wrcell13_mux==1?sd1_d3_io:
			pwm0_pwm_io;

      rule assign_wrsd0_d3_in_on_cell13(wrcell13_mux==0);
        wrsd0_d3_in<=cell13_mux_in;
      endrule


      rule assign_wrsd1_d3_in_on_cell13(wrcell13_mux==1);
        wrsd1_d3_in<=cell13_mux_in;
      endrule

      cell4_mux_out=uart1_tx_io;
      cell5_mux_out=uart1_rx_io;
      cell6_mux_out=twi1_sda_io;
      cell7_mux_out=twi1_scl_io;
      cell14_mux_out=jtag0_tclk_io;
      cell15_mux_out=jtag0_tdo_io;
      cell16_mux_out=jtag0_tdi_io;
      cell17_mux_out=jtag0_tms_io;
      cell18_mux_out=jtag0_tdo_io;

      /*============================================================*/

    interface mux_lines = interface MuxSelectionLines

      method Action  cell0_mux(Bit#(2) in);
         wrcell0_mux<=in;
      endmethod

      method Action  cell1_mux(Bit#(2) in);
         wrcell1_mux<=in;
      endmethod

      method Action  cell2_mux(Bit#(2) in);
         wrcell2_mux<=in;
      endmethod

      method Action  cell3_mux(Bit#(2) in);
         wrcell3_mux<=in;
      endmethod

      method Action  cell8_mux(Bit#(2) in);
         wrcell8_mux<=in;
      endmethod

      method Action  cell9_mux(Bit#(2) in);
         wrcell9_mux<=in;
      endmethod

      method Action  cell10_mux(Bit#(2) in);
         wrcell10_mux<=in;
      endmethod

      method Action  cell11_mux(Bit#(2) in);
         wrcell11_mux<=in;
      endmethod

      method Action  cell12_mux(Bit#(2) in);
         wrcell12_mux<=in;
      endmethod

      method Action  cell13_mux(Bit#(2) in);
         wrcell13_mux<=in;
      endmethod

    endinterface;
    interface peripheral_side = interface PeripheralSide

      method io0_cell=cell0_mux_out;
      method Action  io0_inputval(Bit#(1) in);
         cell0_mux_in<=in;
      endmethod

      method io1_cell=cell1_mux_out;
      method Action  io1_inputval(Bit#(1) in);
         cell1_mux_in<=in;
      endmethod

      method io2_cell=cell2_mux_out;
      method Action  io2_inputval(Bit#(1) in);
         cell2_mux_in<=in;
      endmethod

      method io3_cell=cell3_mux_out;
      method Action  io3_inputval(Bit#(1) in);
         cell3_mux_in<=in;
      endmethod

      method io4_cell=cell4_mux_out;
      method Action  io4_inputval(Bit#(1) in);
         cell4_mux_in<=in;
      endmethod

      method io5_cell=cell5_mux_out;
      method Action  io5_inputval(Bit#(1) in);
         cell5_mux_in<=in;
      endmethod

      method io6_cell=cell6_mux_out;
      method Action  io6_inputval(Bit#(1) in);
         cell6_mux_in<=in;
      endmethod

      method io7_cell=cell7_mux_out;
      method Action  io7_inputval(Bit#(1) in);
         cell7_mux_in<=in;
      endmethod

      method io8_cell=cell8_mux_out;
      method Action  io8_inputval(Bit#(1) in);
         cell8_mux_in<=in;
      endmethod

      method io9_cell=cell9_mux_out;
      method Action  io9_inputval(Bit#(1) in);
         cell9_mux_in<=in;
      endmethod

      method io10_cell=cell10_mux_out;
      method Action  io10_inputval(Bit#(1) in);
         cell10_mux_in<=in;
      endmethod

      method io11_cell=cell11_mux_out;
      method Action  io11_inputval(Bit#(1) in);
         cell11_mux_in<=in;
      endmethod

      method io12_cell=cell12_mux_out;
      method Action  io12_inputval(Bit#(1) in);
         cell12_mux_in<=in;
      endmethod

      method io13_cell=cell13_mux_out;
      method Action  io13_inputval(Bit#(1) in);
         cell13_mux_in<=in;
      endmethod

      method io14_cell=cell14_mux_out;
      method Action  io14_inputval(Bit#(1) in);
         cell14_mux_in<=in;
      endmethod

      method io15_cell=cell15_mux_out;
      method Action  io15_inputval(Bit#(1) in);
         cell15_mux_in<=in;
      endmethod

      method io16_cell=cell16_mux_out;
      method Action  io16_inputval(Bit#(1) in);
         cell16_mux_in<=in;
      endmethod

      method io17_cell=cell17_mux_out;
      method Action  io17_inputval(Bit#(1) in);
         cell17_mux_in<=in;
      endmethod

      method io18_cell=cell18_mux_out;
      method Action  io18_inputval(Bit#(1) in);
         cell18_mux_in<=in;
      endmethod

      method uart0_rx=wruart0_rx;
      method Action  uart0_tx(Bit#(1) in);
         wruart0_tx<=in;
      endmethod

      method uart1_rx=wruart1_rx;
      method Action  uart1_tx(Bit#(1) in);
         wruart1_tx<=in;
      endmethod

      method uart2_rx=wruart2_rx;
      method Action  uart2_tx(Bit#(1) in);
         wruart2_tx<=in;
      endmethod

      method uart3_rx=wruart3_rx;
      method Action  uart3_tx(Bit#(1) in);
         wruart3_tx<=in;
      endmethod

      method Action  spi_sclk(Bit#(1) in);
         wrspi_sclk<=in;
      endmethod
      method Action  spi_mosi(Bit#(1) in);
         wrspi_mosi<=in;
      endmethod
      method Action  spi_ss(Bit#(1) in);
         wrspi_ss<=in;
      endmethod
      method spi_miso=wrspi_miso;

      method Action  twi0_sda_out(Bit#(1) in);
         wrtwi0_sda_out<=in;
      endmethod
      method Action  twi0_sda_outen(Bit#(1) in);
         wrtwi0_sda_outen<=in;
      endmethod
      method twi0_sda_in=wrtwi0_sda_in;
      method Action  twi0_scl_out(Bit#(1) in);
         wrtwi0_scl_out<=in;
      endmethod
      method Action  twi0_scl_outen(Bit#(1) in);
         wrtwi0_scl_outen<=in;
      endmethod
      method twi0_scl_in=wrtwi0_scl_in;

      method Action  twi1_sda_out(Bit#(1) in);
         wrtwi1_sda_out<=in;
      endmethod
      method Action  twi1_sda_outen(Bit#(1) in);
         wrtwi1_sda_outen<=in;
      endmethod
      method twi1_sda_in=wrtwi1_sda_in;
      method Action  twi1_scl_out(Bit#(1) in);
         wrtwi1_scl_out<=in;
      endmethod
      method Action  twi1_scl_outen(Bit#(1) in);
         wrtwi1_scl_outen<=in;
      endmethod
      method twi1_scl_in=wrtwi1_scl_in;

      method Action  sd0_clk(Bit#(1) in);
         wrsd0_clk<=in;
      endmethod
      method Action  sd0_cmd(Bit#(1) in);
         wrsd0_cmd<=in;
      endmethod
      method Action  sd0_d0_out(Bit#(1) in);
         wrsd0_d0_out<=in;
      endmethod
      method Action  sd0_d0_outen(Bit#(1) in);
         wrsd0_d0_outen<=in;
      endmethod
      method sd0_d0_in=wrsd0_d0_in;
      method Action  sd0_d1_out(Bit#(1) in);
         wrsd0_d1_out<=in;
      endmethod
      method Action  sd0_d1_outen(Bit#(1) in);
         wrsd0_d1_outen<=in;
      endmethod
      method sd0_d1_in=wrsd0_d1_in;
      method Action  sd0_d2_out(Bit#(1) in);
         wrsd0_d2_out<=in;
      endmethod
      method Action  sd0_d2_outen(Bit#(1) in);
         wrsd0_d2_outen<=in;
      endmethod
      method sd0_d2_in=wrsd0_d2_in;
      method Action  sd0_d3_out(Bit#(1) in);
         wrsd0_d3_out<=in;
      endmethod
      method Action  sd0_d3_outen(Bit#(1) in);
         wrsd0_d3_outen<=in;
      endmethod
      method sd0_d3_in=wrsd0_d3_in;

      method Action  sd1_clk(Bit#(1) in);
         wrsd1_clk<=in;
      endmethod
      method Action  sd1_cmd(Bit#(1) in);
         wrsd1_cmd<=in;
      endmethod
      method Action  sd1_d0_out(Bit#(1) in);
         wrsd1_d0_out<=in;
      endmethod
      method Action  sd1_d0_outen(Bit#(1) in);
         wrsd1_d0_outen<=in;
      endmethod
      method sd1_d0_in=wrsd1_d0_in;
      method Action  sd1_d1_out(Bit#(1) in);
         wrsd1_d1_out<=in;
      endmethod
      method Action  sd1_d1_outen(Bit#(1) in);
         wrsd1_d1_outen<=in;
      endmethod
      method sd1_d1_in=wrsd1_d1_in;
      method Action  sd1_d2_out(Bit#(1) in);
         wrsd1_d2_out<=in;
      endmethod
      method Action  sd1_d2_outen(Bit#(1) in);
         wrsd1_d2_outen<=in;
      endmethod
      method sd1_d2_in=wrsd1_d2_in;
      method Action  sd1_d3_out(Bit#(1) in);
         wrsd1_d3_out<=in;
      endmethod
      method Action  sd1_d3_outen(Bit#(1) in);
         wrsd1_d3_outen<=in;
      endmethod
      method sd1_d3_in=wrsd1_d3_in;

      method jtag0_tdi=wrjtag0_tdi;
      method jtag0_tms=wrjtag0_tms;
      method jtag0_tclk=wrjtag0_tclk;
      method jtag0_trst=wrjtag0_trst;
      method Action  jtag0_tdo(Bit#(1) in);
         wrjtag0_tdo<=in;
      endmethod

      method jtag1_tdi=wrjtag1_tdi;
      method jtag1_tms=wrjtag1_tms;
      method jtag1_tclk=wrjtag1_tclk;
      method jtag1_trst=wrjtag1_trst;
      method Action  jtag1_tdo(Bit#(1) in);
         wrjtag1_tdo<=in;
      endmethod

      method Action  pwm_pwm(Bit#(1) in);
         wrpwm_pwm<=in;
      endmethod

     endinterface;
   endmodule
endpackage
